library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity PlayerROM is
	port(
		clk_player : in std_logic;
		id_player : in std_logic_vector(3 downto 0);
		x_player : in std_logic_vector(4 downto 0);
		y_player : in std_logic_vector(4 downto 0);
		red_in_player : in std_logic_vector(3 downto 0);
		green_in_player : in std_logic_vector(3 downto 0);
		blue_in_player : in std_logic_vector(3 downto 0);
		red_out_player : out std_logic_vector(3 downto 0);
		green_out_player : out std_logic_vector(3 downto 0);
		blue_out_player : out std_logic_vector(3 downto 0)
	);
end PlayerROM;

architecture PlayerROM_Behav of PlayerROM is

type spriteROM is array(0 to 31) of std_logic_vector(383 downto 0);

constant player1 : spriteROM := (
	x"EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEED97EA8EC9EA8EEEEEEEA8EC9EA8D97EEEEEEEEEEEE730520EEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEE940520EEEEEED97D97EC9EA8D97B76D97EA8EA8EC9D97D97EEEEEE940730730520EEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEE940730520310EEED97EA8EA8D97D97B76D97D97EA8EA8EA8D97EEEEEE940940730730520EEEEEE",
	x"EEEEEEEEEEEEEEEEEE940940730520D97643643EA8643643B76D97643643EA8643643D97EEE940730730520520EEEEEE",
	x"EEEEEEEEEEEEEEE940730730520310D97B76B76EA8B76D97964D97D97B76EA8B76B76D97EEE940940730730520EEEEEE",
	x"EEEEEEEEEEEEEEE940940730730520B76900900900900D97964B76D97900900900900B76B76EEE940520730520EEEEEE",
	x"EEEEEEEEEEEEEEE940730940730520700700700700700700964B76700700700700700700B76EEE940730730520EEEEEE",
	x"EEEEEEEEEEEEEEE940730730520520700CCC700700CCC700643964700CCC700700CCC700B76964730730520EEEEEEEEE",
	x"EEEEEEEEEEEEB76940940730520643B76B76B76B76B76B76643643B76B76B76B76B76B76643964940730520EEEEEEEEE",
	x"EEEEEEEEEB76D97B76940730730B76643643643643643643B76B76643643643643643643B76964940730520EEEEEEEEE",
	x"EEEEEEB76D97964B76940730520643964964B76D97D97B76B76B76B76D97D97B76B76643643B76940730520964EEEEEE",
	x"EEEEEED97B76B76643730730520EEE643964D97B76B76B76964B76D97B76B76964964643EEE940730520B76B76EEEEEE",
	x"EEEB76D97B76643940730520520EEE964643B76B76B76B76964B76B76B76B76964643EEEEEE940730520D97964EEEEEE",
	x"EEE964B76B76964940730730EEEEEE964B76964964964964B76B76964964964643964EEEEEE940730520D97964EEEEEE",
	x"EEE643B76D97B76940730520EEE643964B76D97D97D97D97D97B76B76B76B76964964000EEEEEE730520B76964EEEEEE",
	x"EEEEEE643D97B76B76730520EEE643964B76D97D97D97D97D97D97D97B76B76964964000000EEE730520B76643EEEEEE",
	x"EEEEEEEEE964D97B76D97D97EEE300964B76B76D97D97D97D97D97B76B76B76B76964000000964730520B76643EEEEEE",
	x"EEEEEEEEEEEE643B76B76B76EEE300500964964B76B76B76B76B76B76B76964964300000964D97B76B76964000EEEEEE",
	x"EEEEEEEEEEEEEEE643964964EEE960500500643964964964222964964964643300300000643B76B76B76643000EEEEEE",
	x"EEEEEEEEEEEEEEE730520EEEEEE960B80500500710710643643643643500500300960000000643643643000000EEEEEE",
	x"EEEEEEEEEEEEEEE520EEEEEE530960750B80500710710710710710710500500B80530960000000000000000000EEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEEEEE960B80B80750D90960D90710710710710960B80B80960960000000000000000000EEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEE530960750643B80960D90960D90960D90960D90B80750B80530000000000000000000EEEEEE",
	x"EEEEEEEEEEEEEEEEEE960960960B80643B80D90643D90D90D90D90D90643B80B80643960000000000000000EEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEE960643B80960D90960643960D90643960D90643750B80964000000000000000000EEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEEEEE643B76964960964643643960000D90643964B76B80D97B76000000000000EEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEEEEE643D97D97D90964643000000000D90643964B76B76D97964000000000000EEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEE643964B76B76964643000000000EEEEEE643964B76964964000000000000EEEEEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEE643964964964964643000000EEEEEEEEEEEE643964B76B76000000000000EEEEEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEE964B76B76B76964000000EEEEEEEEEEEEEEE643964964D97D97B76000EEEEEEEEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEE964964964643643000EEEEEEEEEEEEEEE000643643964964964964000EEEEEEEEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEE000000000000000000000EEEEEEEEEEEEEEE000000000000000000000EEEEEEEEEEEEEEEEEEEEE"
);

constant player2 : spriteROM := (
	x"EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEB00D00900EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE00EEEEEEB00E00D00B00900EEEEEEE00EEEEEEEEEEEEEEEEEEEEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE00B00E00D00B00B00900700E00EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEEEEEEEEE00EEEEEEEEEB00200D00B00B00200700EEEEEEE00EEEEEEEEEEEEEEEEEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE00E00E00700200EE0200EE0200500E00E00EEEEEEEEEEEEEEEEEEEEEE00EEEEEE",
	x"EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE700D0020020020090050000B00B00B900900EEEEEEEEEEEEE00EEEEEE",
	x"EEEEEEEEEEEEE00EEEEEEEEEEEEEEE00B00B00E700D00B00200D0090050000E00EB00B00E00E00900EEEE00EEEEEEEEE",
	x"EEEEEEEEEEEEE00EEEEEEEEE900B00B0000E00E00BD00B00200D0090000B00E900900900B00B00E00900EEEEEEEEEEEE",
	x"EEEEEEEEEEEEEEEE00EEE900E00E00B00900B9300E00E00B70000B00E00EB00B93900900ED5C94B00B00900EEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEE900E00B00900900B93B00D00E0000B00B00BB00B00B00B00EB3ED5ED5C94972B00900EEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEE900B00B00900900B93B00D00E00D00D00B00B00B00900900C94EB3ED5EB3972900900EEEEEEEEE",
	x"EEEEEEEEEEEEEEEEEE900B00B00900EB3B00B00000000000E00D00000000000700C94ED5EB3ED5B9397200E00BEEEEEE",
	x"EEEEEEEEEEEEEEEEEEB93EB3EB3EB3200200B00000000000E00D00000000000C94C94EB3EB3ED5C9497200E00BEEEEEE",
	x"EEEEEEEEEEEEEEE00B00E200200200200003B00B00000000E00D00000000700C94C94C94EB3ED5C9497200E00BEEEEEE",
	x"EEEEEEEEEEEEEEE00B00EEB3B93200200003003900B00E00000D00B00900700972B93B93EB3EB3ED5B9397200EEEEEEE",
	x"EEEEEEEEEEEEEEE00BB00E00B00761200003003003B00D00000000900700700761972B93C94EB3ED5C9497200EEEEEEE",
	x"EEEEEEEEEEEEEEE00BB00E00900500003003003999900B00000000700700500500761972B93C94ED5C9497200EEEEEEE",
	x"EEEEEEEEEEEE00EB00E00B00500003003003999999900B00900700700500200999761972B93C94EB3ED597200EEEEEEE",
	x"EEEEEEEEEEEE00EB00E00900500003003003999300300900900700500000200999999761972B93EB3ED597200EEEEEEE",
	x"EEEEEEEEEEEEE00E00900500003003003003999300300999000003999200200200999761972B93C94ED5C94972EEEEEE",
	x"EEEEEEEEE00BB00E00500003003003003300300300999999000003999999200200999100761972B93EB3ED5972EEEEEE",
	x"EEEEEEEEE00B700500500003003003003300300300999000003003003999200000100500761972B93C94ED5972000EEE",
	x"EEEEEEEEE00B00E00E00B003003003003300300300999000003003003999500900900E00003761972C94C94972000EEE",
	x"EEEEEEEEE00B00E00E00B003003003700E00300000000003003003003700700B00E00700003003761972C94972000EEE",
	x"EEEEEE00B00B00E00E00E003003003700900700900500003003003003003500900E00700003003003761972972000EEE",
	x"EEEEEE00B00B00E00B003003003003700900700900500003003003003003500B00E00700003003003003972972000EEE",
	x"EEEEEE00B00E00E00B003003003003003700E00900500003003003003003500900E00700003003003003761761000EEE",
	x"EEE00B00B00E00E00B003003003003003700E00700500003003003000000500700900B00E00000000000000761EEEEEE",
	x"EEE00B00B00E00E00B003000000000000900900700500003003000000000000500700900B00E00000000EEEEEEEEEEEE",
	x"EEE00B00B00E00E00B000000000000700E00900500500000000000000000000000000700700700000EEEEEEEEEEEEEEE",
	x"EEEEEE00B00E00E00B000000000000700E00500500000000000000000EEEEEEEEE000000000000EEEEEEEEEEEEEEEEEE",
	x"EEEEEEEEEEEE000000000000000000900900500000000000EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE"
);

begin
	player_proc : process(clk_player)
	
	variable x_int : integer range 0 to 31 := 0;
	variable y_int : integer range 0 to 31 := 0;
	variable sprite_idx : integer range 0 to 383 := 0;
	variable red : std_logic_vector(3 downto 0) := x"0";
	variable green : std_logic_vector(3 downto 0) := x"0";
	variable blue : std_logic_vector(3 downto 0) := x"0";
	
	begin
		if(clk_player'event and clk_player = '1') then
			x_int := to_integer(unsigned(x_player));
			y_int := to_integer(unsigned(y_player));
			sprite_idx := 383 - 6 * x_int;
			case id_player is
				when x"2" => 
					red := player1(y_int)(sprite_idx downto (sprite_idx - 3));
					green := player1(y_int)((sprite_idx - 4) downto (sprite_idx - 7));
					blue := player1(y_int)((sprite_idx - 8) downto (sprite_idx - 11));
				when x"3" =>
					red := player2(y_int)(sprite_idx downto (sprite_idx - 3));
					green := player2(y_int)((sprite_idx - 4) downto (sprite_idx - 7));
					blue := player2(y_int)((sprite_idx - 8) downto (sprite_idx - 11));
				when others =>
					red := x"E";
					green := x"E";
					blue := x"E";
			end case;
			
			if(red = x"E" and green = x"E" and blue = x"E") then
				red_out_player <= red_in_player;
				green_out_player <= green_in_player;
				blue_out_player <= blue_in_player;
			else
				red_out_player <= red;
				green_out_player <= green;
				blue_out_player <= blue;
			end if;
		end if;
	end process player_proc;


end PlayerROM_Behav;

